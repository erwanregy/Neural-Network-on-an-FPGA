`include "include.svh"

module test_rom;

    // ROM

    localparam int NUM_WEIGHTS = 784;
    localparam string WEIGHTS_FILE = "weights.mem";

    logic clock, reset;
    logic [$clog2(NUM_WEIGHTS)-1:0] weight_num;
    logic signed [INT_WIDTH-1:-FRAC_WIDTH] weight;

    rom #(
        .WIDTH(INT_WIDTH + FRAC_WIDTH),
        .DEPTH(NUM_WEIGHTS),
        .FILE(WEIGHTS_FILE)
    ) parameters (
        .clock(clock),
        .address(weight_num),
        .out(weight)
    );


    // Clock generator

    clock_generator cg (.*);


    // Testbench

    initial begin
        #RESET_PERIOD;
        for (int i = 0; i < NUM_WEIGHTS; i++) begin
            weight_num = i;
            #CLOCK_PERIOD;
        end
        $finish;
    end

endmodule